module decoder_2x4(input en,input [1:0]a,output reg [3:0]y);

always@ (en or a)begin

if (en == 0)
y=4'b0000;
else begin
case(a)
      2'b00:y=4'b0001;
      2'b01:y=4'b0010;
      2'b10:y=4'b0100;
      2'b11:y=4'b1000;
default:y[3:0]=4'b0000;
endcase
end
end
endmodule
