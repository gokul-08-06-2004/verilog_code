module half_sub(input a,b,output diff,barrow);

assign {barrow,diff}=a-b;

endmodule

