//48. Use $dumpfile and $dumpvars to generate waveform for a NOT gate.

module not_gate(input a,output y);

assign y=~a;
endmodule
