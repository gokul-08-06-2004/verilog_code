module inverter_tb;
reg a;                                                                                                                  output y;                                                                                                               inverter dut(a,y);                                                                                                                                                                                                                              initial begin                                                                                                                                                                                                                                   $monitor("a=%b",y);                                                                                                                                                                                                                             a=0;                                                                                                                    a=1;                                                                                                                                                                                                                                            $finish;                                                                                                                end                                                                                                                     endmodule          
