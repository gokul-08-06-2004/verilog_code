module basic_gates(input a,b, output y);
nor (y,a,b);
endmodule
