module encoder_tb;
reg [7:0]a;
wire [2:0]y;

encoder_8x1 dut(a,y);

initial begin

$monitor("a[7]=%b a[6]=%b a[5]=%b a[4]=%b a[3]=%b a[2]=%b a[1]=%b a[0]=%b | y[2]=%b y[1]=%b y[0]=%b",a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],y[2],y[1],y[0]);
$dumpfile("encoder.vcd");
$dumpvars();

a[7]=0; a[6]=0; a[5]=0; a[4]=0; a[3]=0; a[2]=0; a[1]=0; a[0]=1; #10
a[7]=0; a[6]=0; a[5]=0; a[4]=0; a[3]=0; a[2]=0; a[1]=1; a[0]=0; #10
a[7]=0; a[6]=0; a[5]=0; a[4]=0; a[3]=0; a[2]=1; a[1]=0; a[0]=0; #10
a[7]=0; a[6]=0; a[5]=0; a[4]=0; a[3]=1; a[2]=0; a[1]=0; a[0]=0; #10
a[7]=0; a[6]=0; a[5]=0; a[4]=1; a[3]=0; a[2]=0; a[1]=0; a[0]=0; #10
a[7]=0; a[6]=0; a[5]=1; a[4]=0; a[3]=0; a[2]=0; a[1]=0; a[0]=0; #10
a[7]=0; a[6]=1; a[5]=0; a[4]=0; a[3]=0; a[2]=0; a[1]=0; a[0]=0; #10
a[7]=1; a[6]=0; a[5]=0; a[4]=0; a[3]=0; a[2]=0; a[1]=0; a[0]=0; #10

$finish;
end 
endmodule

