//14. Create a pipelined register using non-blocking assignments.

module pipelined()
