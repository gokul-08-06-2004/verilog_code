
module basic_gates(input a,b, output y);
nand (y,a,b);
endmodule
