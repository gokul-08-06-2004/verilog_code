module mux_8x1_tb();

reg i0,i1,i2,i3,i4,i5,i6,i7,s0,s1,s2;
wire y;

mux_8x1 dut(i0,i1,i2,i3,i4,i5,i6,i7,s0,s1,s2,y);

initial begin 

$monitor("i0=%b i1=%b i2=%b i3=%b i4=%b i5=%b i6=%b i7=%b s0=%b s1=%b s2=%b y=%b ",i0,i1,i2,i3,i4,i5,i6,i7,s0,s1,s2,y);
$dumpfile("mux_8x1.vcd");
$dumpvars();

i0=1; i1=1; i2=1; i3=0; i4=1; i5=0; i6=1; i7=1;

s0=0; s1=0; s2=0; #10
s0=0; s1=0; s2=1; #10
s0=0; s1=1; s2=0; #10
s0=0; s1=1; s2=1; #10
s0=1; s1=0; s2=0; #10
s0=1; s1=0; s2=1; #10
s0=1; s1=1; s2=0; #10
s0=1; s1=1; s2=1; #10


$finish;
end 
endmodule 
