module add_tb;
reg a,b;
wire out;

add dut(a,b,out);

initial begin
$monitor("Time=%0t a=%b b=%b out=%b ",$time, a,b,out);

a=0; b=0;#10
a=0; b=1;#10
a=1; b=0; #10
a=1; b=1; #10

$finish;
end
endmodule
