//1. Write a Verilog module using a continuous assignment to implement out = a & b.

module conti(input a,b,output out);

assign out= a&b;

endmodule
