module int();
integer b;
initial begin
b=-'d12/3;#10
$finish;
end
endmodule
