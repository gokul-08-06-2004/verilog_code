module basic_gates_tb;

reg a,b;
wire y;

basic_gates dut(a,b,y);

initial begin

$monitor("a=%b | b=%b y=%b",a,b,y);
$dumpfile("basic_gates.vcd");
$dumpvars();


a=0; b=0; #10
a=0; b=1; #10
a=1; b=0; #10
a=1; b=1; #10

$finish;
end
endmodule
