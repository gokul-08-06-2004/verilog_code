//51. Write a testbench for a 1-bit NOT gate.

module not_gate(input a,output y);

assign y=~a;

endmodule
