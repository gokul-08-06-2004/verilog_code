module encoder(input [3:0]a,output [1:0]y);

assign y[1:0]=(a==4'b0001)?2'b00:
              (a==4'b0010)?2'b01:
              (a==4'b0100)?2'b10:
                           2'b11;

endmodule
